// hazard.v

// This module determines if pipeline stalls or flushing are required

// TODO: declare propoer input and output ports and implement the
// hazard detection unit

module hazard ( //UNDONE
    input [4:0] rs1_id,
    input [4:0] rs2_id,
    input [4:0] rd_ex,

    output flush, stall
);


endmodule
